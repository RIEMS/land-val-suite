netcdf init {
dimensions:
	west_east = 1 ;
	south_north = 1 ;
	soil_layers = 4 ;
	snow_layers = 3 ;
variables:
	double XLAT(south_north, west_east) ;
		XLAT:long_name = "latitude" ;
		XLAT:units = "degree_north" ;
		XLAT:standard_name = "latitude" ;
	double XLONG(south_north, west_east) ;
		XLONG:long_name = "longitude" ;
		XLONG:units = "degree_east" ;
		XLONG:standard_name = "longitude" ;
	byte XLAND(south_north, west_east) ;
		XLAND:long_name = "land sea mask" ;
		XLAND:units = "-" ;
		XLAND:standard_name = "land_binary_mask" ;
		XLAND:_FillValue = 0b ;
		XLAND:valid_range = 1b, 2b ;
		XLAND:flag_value = 1b, 2b ;
		XLAND:flag_meanings = "land sea" ;
	float CANLIQ(south_north, west_east) ;
		CANLIQ:long_name = "canopy_liquid_water_amount" ;
		CANLIQ:units = "kg m-2" ;
		CANLIQ:_FillValue = NaN ;
	float CANICE(south_north, west_east) ;
		CANICE:standard_name = "canopy_snow_amount" ;
		CANICE:units = "kg m-2" ;
		CANICE:_FillValue = NaN ;
	float TV(south_north, west_east) ;
		TV:standard_name = "canopy_temperature" ;
		TV:units = "K" ;
		TV:_FillValue = NaN ;
	float TG(south_north, west_east) ;
		TG:standard_name = "surface_temperature" ;
		TG:units = "K" ;
		TG:_FillValue = NaN ;
	int NSNOW(south_north, west_east) ;
		NSNOW:long_name = "snow_layer_count" ;
		NSNOW:units = "1" ;
		NSNOW:_FillValue = -1 ;
	float SNOW(south_north, west_east) ;
		SNOW:standard_name = "surface_snow_amount" ;
		SNOW:units = "kg m-2" ;
		SNOW:_FillValue = NaN ;
	float SNOWH(south_north, west_east) ;
		SNOWH:standard_name = "surface_snow_thickness" ;
		SNOWH:units = "m" ;
		SNOWH:_FillValue = NaN ;
	float DZSNOW(snow_layers, south_north, west_east) ;
		DZSNOW:standard_name = "surface_snow_thickness" ;
		DZSNOW:units = "m" ;
		DZSNOW:_FillValue = NaN ;
	float SNOWT(snow_layers, south_north, west_east) ;
		SNOWT:standard_name = "snow_temperature" ;
		SNOWT:units = "K" ;
		SNOWT:_FillValue = NaN ;
	float SNOWLIQ(snow_layers, south_north, west_east) ;
		SNOWLIQ:standard_name = "liquid_water_content_of_surface_snow" ;
		SNOWLIQ:units = "kg m-2" ;
		SNOWLIQ:_FillValue = NaN ;
	float SNOWICE(snow_layers, south_north, west_east) ;
		SNOWICE:standard_name = "solid_water_content_of_surface_snow" ;
		SNOWICE:units = "kg m-2" ;
		SNOWICE:_FillValue = NaN ;
	float SOILT(soil_layers, south_north, west_east) ;
		SOILT:long_name = "soil layer temperature" ;
		SOILT:units = "K" ;
		SOILT:_FillValue = NaN ;
	float SOILM(soil_layers, south_north, west_east) ;
		SOILM:long_name = "soil layer moisture content" ;
		SOILM:units = "m3 m-3" ;
		SOILM:_FillValue = NaN ;
		SOILM:valid_range = 0., 1. ;
	float SOILMLIQ(soil_layers, south_north, west_east) ;
		SOILMLIQ:long_name = "soil layer moisture liquid content" ;
		SOILMLIQ:units = "m3 m-3" ;
		SOILMLIQ:_FillValue = NaN ;
		SOILMLIQ:valid_range = 0., 1. ;
	float WA(south_north, west_east) ;
		WA:long_name = "groundwater_amount" ;
		WA:units = "kg m-2" ;
		WA:_FillValue = NaN ;
	float WT(south_north, west_east) ;
		WT:long_name = "water_storage_in_saturated_soil_and_groundwater" ;
		WT:units = "kg m-2" ;
		WT:_FillValue = NaN ;
	float ZWT(south_north, west_east) ;
		ZWT:long_name = "water_table_depth" ;
		ZWT:units = "m" ;
		ZWT:_FillValue = NaN ;
	float LAI(south_north, west_east) ;
		LAI:long_name = "leaf area index" ;
		LAI:units = "m2 m-2" ;
		LAI:standard_name = "leaf_area_index" ;
		LAI:_FillValue = NaN ;
	float SAI(south_north, west_east) ;
		SAI:long_name = "stem area index" ;
		SAI:units = "m2 m-2" ;
		SAI:standard_name = "stem_area_index" ;
		SAI:_FillValue = NaN ;
	float LFMASS(south_north, west_east) ;
		LFMASS:long_name = "leaf_mass" ;
		LFMASS:units = "g m-2" ;
		LFMASS:_FillValue = NaN ;
	float RTMASS(south_north, west_east) ;
		RTMASS:long_name = "root_mass" ;
		RTMASS:units = "g m-2" ;
		RTMASS:_FillValue = NaN ;
	float STMASS(south_north, west_east) ;
		STMASS:long_name = "stem_mass" ;
		STMASS:units = "g m-2" ;
		STMASS:_FillValue = NaN ;
	float WDMASS(south_north, west_east) ;
		WDMASS:long_name = "wood_mass" ;
		WDMASS:units = "g m-2" ;
		WDMASS:_FillValue = NaN ;
	float STBLCP(south_north, west_east) ;
		STBLCP:long_name = "stable_carbon_pool" ;
		STBLCP:units = "g m-2" ;
		STBLCP:_FillValue = NaN ;
	float FASTCP(south_north, west_east) ;
		FASTCP:long_name = "fast_carbon_pool" ;
		FASTCP:units = "g m-2" ;
		FASTCP:_FillValue = NaN ;

// global attributes:
		:title = "Bondville surface meteorological data" ;
data:

 XLAT =
  40.01 ;

 XLONG =
  -88.37 ;

 CANLIQ =
  0.01 ;

 CANICE =
  0.00 ;

 TV =
  263.7 ;

 TG =
  263.7 ;

 NSNOW =
  0 ;

 SNOW =
  1 ;

 SNOWH =
  0.01 ;

 DZSNOW =
  0.01,
  0.00,
  0.00 ;

 SNOWT =
  273.15,
  273.15,
  273.15 ;

 SNOWLIQ =
  0.00,
  0.00,
  0.00 ;

 SNOWICE =
  1.0,
  0.00,
  0.00 ;

 SOILT =
  266.1,
  274,
  276.9,
  279.9 ;

 SOILM =
  0.298,
  0.294,
  0.271,
  0.307 ;

 SOILMLIQ =
  0.298,
  0.294,
  0.271,
  0.307 ;

 WA =
  4900.0 ;

 WT =
  4900.0 ;

 ZWT =
  2.5 ;

 LAI =
  2 ;

 SAI =
  0.2 ;

 LFMASS =
  0.83 ;

 STMASS =
  16.67 ;

 RTMASS =
  500.0 ;

 WDMASS =
  500.0 ;

 STBLCP =
  1000.0 ;

 FASTCP =
  1000.0 ;
}
